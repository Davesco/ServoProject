--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   23:02:29 09/25/2012
-- Design Name:   
-- Module Name:   C:/Users/Administrador/Desktop/Lab_electroII/uart/uart/Tb1_Rx.vhd
-- Project Name:  uart
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: RX_module
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Tb1_Rx IS
END Tb1_Rx;
 
ARCHITECTURE behavior OF Tb1_Rx IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT RX_module
    PORT(
         clk : IN  std_logic;
         serie : IN  std_logic;
         
			encb : out  STD_LOGIC;
         data : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal serie : std_logic := '0';

 	--Outputs
   signal data : std_logic_vector(7 downto 0);
	signal encb : STD_LOGIC;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: RX_module PORT MAP (
          clk => clk,
          serie => serie,
          data => data,
			 encb => encb 
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
			serie<='1';
		wait for 10 ns;	
			serie<='1';
		wait for 10 ns;	
			serie<='1';
		wait for 10 ns;	
			serie<='1';
		wait for 10 ns;	
			serie<='0';
		wait for 10 ns;	
			serie<='1';
		wait for 10 ns;	
			serie<='0';
		wait for 10 ns;
			serie<='1';
		wait for 10 ns;
			serie<='1';
		wait for 10 ns;
			serie<='0';
		wait for 10 ns;
			serie<='1';
		wait for 10 ns;
			serie<='1';
		wait for 10 ns;
			serie<='0';
		wait for 10 ns;
			serie<='1';
		wait for 10 ns;	
			serie<='1';	
wait for 5 ns;		
		

      -- insert stimulus here 

      wait;
   end process;

END;
